/*------------------------------------------------------------------------------
 * File          : main.sv
 * Project       : RTL
 * Author        : epebar
 * Creation date : Jan 20, 2023
 * Description   :
 *------------------------------------------------------------------------------*/

module main #(
	parameter WINDOW_SIZE              = 128,
	          KMER_SIZE                = 16,
	          SKETCH_SIZE              = 16,
	          NUM_OF_BUCKETS           = 256,
	          BUCKET_SIZE              = 16,
	          MAX_WINDOWS_IN_REFERENCE = 512,
	          MAX_WINDOWS_IN_READ      = 16,
	          WINDOWS_PER_QUERY        = 1 // For dealing with multiple read windows at once using posible future query module
) ();


// Wires
// ==================================================
// Interface between main and top level
logic                            hashing_is_done;
logic                            calculate_matched_window;
logic                            reset_stats;
logic                            clk;
logic                            reset_hash_table;
logic  [1:0]                     window       [0:WINDOW_SIZE-1]; // consists of WINDOW_SIZE kmers
logic  [31:0]                    window_id;
logic                        	 ready_for_hashing;
logic                        	 reset_window_hasher;
logic                            is_insert;
logic                            is_query;
logic signed [31:0]              matched_window_id;
// ==================================================


// Top Level Instantiation
// ==================================================
top_level top_level_inst (
	.calculate_matched_window(calculate_matched_window),
	.reset_stats(reset_stats),
	.clk(clk),
	.reset_hash_table(reset_hash_table),
	.window(window),
	.window_id(window_id),
	.ready_for_hashing(ready_for_hashing),
	.reset_window_hasher(reset_window_hasher),
	.is_insert(is_insert),
	.is_query(is_query),
	
	.hashing_is_done(hashing_is_done),
	.matched_window_id(matched_window_id)
);
defparam top_level_inst.WINDOW_SIZE = WINDOW_SIZE;
defparam top_level_inst.KMER_SIZE = KMER_SIZE;
defparam top_level_inst.SKETCH_SIZE = SKETCH_SIZE;
defparam top_level_inst.NUM_OF_BUCKETS = NUM_OF_BUCKETS;
defparam top_level_inst.BUCKET_SIZE = BUCKET_SIZE;
defparam top_level_inst.MAX_WINDOWS_IN_REFERENCE = MAX_WINDOWS_IN_REFERENCE;
defparam top_level_inst.MAX_WINDOWS_IN_READ = MAX_WINDOWS_IN_READ;
defparam top_level_inst.WINDOWS_PER_QUERY = WINDOWS_PER_QUERY;
// ==================================================


always #1 clk=~clk; // Creation of a clock


task reset_all();
	clk = 1'b0;
	
	reset_hash_table = 1'b1;
	reset_window_hasher = 1'b1;
	reset_stats = 1'b1;
	
	calculate_matched_window = 1'b0;
	window = '{default: '0};
	window_id = 0;
	ready_for_hashing = 1'b0;
	is_insert = 1'b0;
	is_query = 1'b0;
	
	#4;
	
	reset_hash_table = 1'b0;
	reset_window_hasher = 1'b0;
	reset_stats = 1'b0;
endtask


// Variables
// ==================================================
int char;
int fd;
int read_file_number;
int fseek_output;
logic was_reading_cancelled;

string read_file_name;
// ==================================================


// Reads windows from given reference or read file and feed them to hardware
task read_and_feed_windows(int fd, logic is_reference);
	
	window_id = 0; // Current window index
	was_reading_cancelled = 1'b0;
	
	reset_window_hasher = 1'b1;
	reset_stats = 1'b1;
	#4;
	reset_window_hasher = 1'b0;
	reset_stats = 1'b0;
	
	while (1'b1) begin
		
		// Assign to window according to nucleotides in file
		// $display("Beginning reading window #%0d...", window_id); // TODO: This is a debugging print
		for (int j = 0; j < WINDOW_SIZE && !was_reading_cancelled; j++) begin
			
			char = $fgetc(fd);
			case (char)
				"A": window[j] = 2'b00;
				"C": window[j] = 2'b01;
				"G": window[j] = 2'b10;
				"T": window[j] = 2'b11;
				default: begin
					// $display("Ignoring reading of window #%0d. It's too short.", window_id);  // TODO: This is a debugging print
					was_reading_cancelled = 1'b1;
				end
			endcase
		end
		
		// To solve eof final chars (like char 10):
		char = $fgetc(fd);
		char = $fgetc(fd);
		
		
		if (!was_reading_cancelled) begin
			
			// $display("Finished reading window #%0d.", window_id); // TODO: This is a debugging print
			// $display("Beginning hashing..."); // TODO: This is a debugging print
			
			ready_for_hashing = 1'b1;
			wait (hashing_is_done == 1'b1)
			// $display("Hashing is done."); // TODO: This is a debugging print
			ready_for_hashing = 1'b0;
			
			if (is_reference) begin
				
				is_insert = 1'b1;
				#4;
				is_insert = 1'b0;
				#4;
			end
			else begin
				
				is_query = 1'b1;
				#4;
				is_query = 1'b0;
				#4;
			end
		end
		
		if ($feof(fd) || was_reading_cancelled) begin
			
			if (!is_reference) begin
				
				calculate_matched_window = 1'b1;
				#4;
				$display("Finished querying read.");
				if (matched_window_id != -1) begin
					
					$display("Matched window id is: %0d.", matched_window_id);
				end
				else begin
					
					$display("No matching window was found.");
				end
				calculate_matched_window = 1'b0;
			end
			else begin
				
				$display("Finished inserting reference.");
			end
			
			return;
		end
		else begin
			
			window_id++;
			fseek_output = $fseek(fd, (WINDOW_SIZE - KMER_SIZE + 1) * window_id, 0);
			if (fseek_output > 0) begin
				
				$display("fseek error");
				$fclose(fd);
				$finish;
			end

			reset_window_hasher = 1'b1;
			#4;
			reset_window_hasher = 1'b0;
		end
		
	end
endtask


// Main
// ==================================================
initial begin
	reset_all();
	
	// Open and insert reference file
	$display("Beginning to read reference file");
	fd = $fopen("./reference_sv.txt", "r");
	if (fd == 0) begin
		
		$display("Could not open reference_sv");
		$finish;
	end
	read_and_feed_windows(fd, 1'b1);
	$fclose(fd);
	
	// Open and query read files
	read_file_number = 0;
	while (1'b1) begin
		
		$sformat(read_file_name,"./read_files/read_sv_%0d.txt",read_file_number);
		fd = $fopen(read_file_name, "r");
		
		if (fd == 0) begin
			
			$display("Done.");
			$finish;
		end
		
		$display("Beginning to query read file #%0d", read_file_number);	
		read_and_feed_windows(fd, 1'b0);
		$fclose(fd);
		
		read_file_number++;
	end	
end
// ==================================================

endmodule
