/*------------------------------------------------------------------------------
 * File          : window_hasher.sv
 * Project       : RTL
 * Author        : epebar
 * Creation date : Nov 29, 2022
 * Description   :
 *------------------------------------------------------------------------------*/

module window_hasher #(
	parameter SKETCH_SIZE         =16,
	          NUM_OF_BUCKETS      =256,
	          WINDOW_SIZE         =128,
	          KMER_SIZE           =16
) (
	input	logic                        clk,
	input	logic                        reset_window_hasher,
	input	logic                        ready_for_hashing,
	input logic  [1:0]                     window        [0:WINDOW_SIZE-1], // consists of WINDOW_SIZE kmers
	
	output logic [$clog2(NUM_OF_BUCKETS)-1:0] hashed_sketch [0:SKETCH_SIZE-1], // vector of SKETCH_SIZE size with each value representing the value of the K-mer after h2 is applied on it
	output logic                           hashing_is_done                  // turns on for one clock cycle when ready
);

logic [31:0] h1_all_kmers  [0:WINDOW_SIZE - KMER_SIZE]; // h1 run on all possible kmers
logic [$clog2(NUM_OF_BUCKETS)-1:0] h2_all_kmers  [0:WINDOW_SIZE - KMER_SIZE]; // h2 run on all possible kmers

logic is_hashing_active;

genvar i;
generate
	for (i = 0 ; i <= WINDOW_SIZE - KMER_SIZE; i++) begin
		hasher u0 (
			.kmer(window[i:i + KMER_SIZE - 1]),
			.h1  (h1_all_kmers[i]            ),
			.h2  (h2_all_kmers[i]            )
		);
	end
endgenerate

logic [31:0] h1_sketch [0:SKETCH_SIZE-1];

logic [31:0] currentSmallest;

logic [31:0] index_in_h1_sketch;
logic [31:0] index_in_h1_all_kmers;

always @(posedge clk or posedge reset_window_hasher) begin
	
	if (reset_window_hasher) begin
		
		currentSmallest = 0;
		index_in_h1_sketch = 0;
		index_in_h1_all_kmers = 0;
		is_hashing_active = 1'b0;
		hashing_is_done = 1'b0;
		hashed_sketch = '{default: '0};
	end
	
	else if (ready_for_hashing == 1'b1 && is_hashing_active == 1'b0) begin
		
		is_hashing_active = 1'b1;
	end
	
	else if (is_hashing_active == 1'b1 && hashing_is_done == 1'b0) begin
		
		if (index_in_h1_all_kmers == 0) begin
			
			h1_sketch[index_in_h1_sketch] = -1;
		end
		
		if (h1_all_kmers[index_in_h1_all_kmers] > currentSmallest
				&& h1_all_kmers[index_in_h1_all_kmers] <= h1_sketch[index_in_h1_sketch]) begin
			
			h1_sketch[index_in_h1_sketch] = h1_all_kmers[index_in_h1_all_kmers];
			hashed_sketch[index_in_h1_sketch] = h2_all_kmers[index_in_h1_all_kmers];
		end
		
		if (index_in_h1_all_kmers == WINDOW_SIZE - KMER_SIZE) begin
			
			if (index_in_h1_sketch == SKETCH_SIZE - 1) begin
				
				hashing_is_done = 1'b1;
			end
			
			else begin
				
				currentSmallest = h1_sketch[index_in_h1_sketch];
				index_in_h1_sketch += 1;
				index_in_h1_all_kmers = 0;
				
			end
		end
		
		else begin
			
			index_in_h1_all_kmers += 1;
		end
	end
end
endmodule
