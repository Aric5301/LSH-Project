/*------------------------------------------------------------------------------
 * File          : hash_table_tb.sv
 * Project       : RTL
 * Author        : epebar
 * Creation date : Sep 24, 2022
 * Description   :
 *------------------------------------------------------------------------------*/

module hash_table_tb #(
	parameter SKETCH_SIZE         =16,
	          NUM_OF_BUCKETS      =256,
	          BUCKET_SIZE         =16,
			  MAX_WINDOWS_IN_REFERENCE = 512
) ();

logic clk;
logic reset_hash_table;
logic is_insert;
logic is_query;
logic [31:0] window_id;
logic [$clog2(NUM_OF_BUCKETS)-1:0] hashed_sketch [0:SKETCH_SIZE-1]; // vector of SKETCH_SIZE size with each value representing the value of the K-mer after h2 is applied on it

logic [31:0] count_bus [0:MAX_WINDOWS_IN_REFERENCE-1]; // currently supports up to 1024 windows

// local parameters, temp as output
logic [31:0] theTable [0:NUM_OF_BUCKETS-1][0:BUCKET_SIZE-1]; // NUM_OF_BUCKETS buckets of BUCKET_SIZE size
logic [31:0] tableLength [0:NUM_OF_BUCKETS-1]; // current length of each bucket

hash_table U1 (.*);

initial begin
	$monitor ("@%g clk= %b reset= %b, isInsert= %b, isQuery= %b, windowID= %d, theTable[0][0]= %d, tableLength[0]= %d, tableLength[1]= %d, countBus[0]= %d, countBus[14]= %d",
			$time,clk,reset_hash_table,is_insert,is_query, window_id, theTable[0][0], tableLength[0], tableLength[1], count_bus[0], count_bus[14]);
	
	
	clk = 1'b0;
	reset_hash_table = 1'b0;
	is_insert = 1'b0;
	is_query = 1'b0;
	window_id = 0;
	
	hashed_sketch[0] = 8'd0;
	hashed_sketch[1] = 8'd0;
	hashed_sketch[2] = 8'd0;
	hashed_sketch[3] = 8'd0;
	hashed_sketch[4] = 8'd0;
	hashed_sketch[5] = 8'd0;
	hashed_sketch[6] = 8'd0;
	hashed_sketch[7] = 8'd0;
	hashed_sketch[8] = 8'd0;
	hashed_sketch[9] = 8'd0;
	hashed_sketch[10] = 8'd0;
	hashed_sketch[11] = 8'd0;
	hashed_sketch[12] = 8'd0;
	hashed_sketch[13] = 8'd0;
	hashed_sketch[14] = 8'd0;
	hashed_sketch[15] = 8'd0;
	
	#2;
	
	reset_hash_table = 1'b1;
	#2;
	reset_hash_table = 1'b0;
	#2;
	window_id = 14;
	is_insert = 1'b1;
	clk = 1'b1;
	#2;
	window_id = 0;
	is_insert = 1'b0;
	clk = 1'b0;
	#2;
	is_query = 1'b1;
	clk = 1'b1;
	#2;
	is_query = 1'b0;
	clk = 1'b0;
	#2;
	
	$finish;
end
endmodule
